`timescale 1ns / 1ps
module datapath_sim(

	reg clock, rst;

    );
endmodule
